module mix_nibbles(cipher,text);
input [63:0]cipher;
output [63:0]text;	

assign text = cipher;
endmodule