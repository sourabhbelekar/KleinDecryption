// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 15.0.0 Build 145 04/22/2015 Patches 0.01we SJ Web Edition"
// CREATED		"Sun Sep 22 15:50:34 2019"

module multi_full_v(
	a,
	b,
	r
);


input wire	[0:7] a;
input wire	[0:7] b;
output wire	[0:7] r;

wire	[0:7] r_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_176;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_110;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_116;
wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_118;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_143;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_145;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_148;
wire	SYNTHESIZED_WIRE_149;
wire	SYNTHESIZED_WIRE_150;
wire	SYNTHESIZED_WIRE_151;
wire	SYNTHESIZED_WIRE_152;
wire	SYNTHESIZED_WIRE_153;
wire	SYNTHESIZED_WIRE_154;
wire	SYNTHESIZED_WIRE_155;
wire	SYNTHESIZED_WIRE_156;
wire	SYNTHESIZED_WIRE_157;
wire	SYNTHESIZED_WIRE_158;
wire	SYNTHESIZED_WIRE_159;
wire	SYNTHESIZED_WIRE_160;
wire	SYNTHESIZED_WIRE_161;
wire	SYNTHESIZED_WIRE_162;
wire	SYNTHESIZED_WIRE_163;
wire	SYNTHESIZED_WIRE_164;
wire	SYNTHESIZED_WIRE_165;
wire	SYNTHESIZED_WIRE_166;
wire	SYNTHESIZED_WIRE_167;
wire	SYNTHESIZED_WIRE_168;
wire	SYNTHESIZED_WIRE_169;
wire	SYNTHESIZED_WIRE_170;
wire	SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_172;
wire	SYNTHESIZED_WIRE_173;
wire	SYNTHESIZED_WIRE_174;
wire	SYNTHESIZED_WIRE_175;

assign	SYNTHESIZED_WIRE_176 = 0;




multiplication_block	b2v_inst(
	.b1(b[0]),
	.b2(b[1]),
	.b3(b[2]),
	.b4(b[3]),
	.b5(b[4]),
	.b6(b[5]),
	.b7(b[6]),
	.b8(b[7]),
	.a1(a[0]),
	.a2(a[1]),
	.a3(a[2]),
	.a4(a[3]),
	.a5(a[4]),
	.a6(a[5]),
	.a7(a[6]),
	.a8(a[7]),
	.r1(SYNTHESIZED_WIRE_176),
	.r2(SYNTHESIZED_WIRE_176),
	.r3(SYNTHESIZED_WIRE_176),
	.r4(SYNTHESIZED_WIRE_176),
	.r5(SYNTHESIZED_WIRE_176),
	.r6(SYNTHESIZED_WIRE_176),
	.r7(SYNTHESIZED_WIRE_176),
	.r8(SYNTHESIZED_WIRE_176),
	.bo_1(SYNTHESIZED_WIRE_8),
	.bo_2(SYNTHESIZED_WIRE_9),
	.bo_3(SYNTHESIZED_WIRE_10),
	.bo_4(SYNTHESIZED_WIRE_11),
	.bo_5(SYNTHESIZED_WIRE_12),
	.bo_6(SYNTHESIZED_WIRE_13),
	.bo_7(SYNTHESIZED_WIRE_14),
	.bo_8(SYNTHESIZED_WIRE_15),
	.ao_1(SYNTHESIZED_WIRE_16),
	.ao_2(SYNTHESIZED_WIRE_17),
	.ao_3(SYNTHESIZED_WIRE_18),
	.ao_4(SYNTHESIZED_WIRE_19),
	.ao_5(SYNTHESIZED_WIRE_20),
	.ao_6(SYNTHESIZED_WIRE_21),
	.ao_7(SYNTHESIZED_WIRE_22),
	.ao_8(SYNTHESIZED_WIRE_23),
	.ro_1(SYNTHESIZED_WIRE_24),
	.ro_2(SYNTHESIZED_WIRE_25),
	.ro_3(SYNTHESIZED_WIRE_26),
	.ro_4(SYNTHESIZED_WIRE_27),
	.ro_5(SYNTHESIZED_WIRE_28),
	.ro_6(SYNTHESIZED_WIRE_29),
	.ro_7(SYNTHESIZED_WIRE_30),
	.ro_8(SYNTHESIZED_WIRE_31));


multiplication_block	b2v_inst1(
	.b1(SYNTHESIZED_WIRE_8),
	.b2(SYNTHESIZED_WIRE_9),
	.b3(SYNTHESIZED_WIRE_10),
	.b4(SYNTHESIZED_WIRE_11),
	.b5(SYNTHESIZED_WIRE_12),
	.b6(SYNTHESIZED_WIRE_13),
	.b7(SYNTHESIZED_WIRE_14),
	.b8(SYNTHESIZED_WIRE_15),
	.a1(SYNTHESIZED_WIRE_16),
	.a2(SYNTHESIZED_WIRE_17),
	.a3(SYNTHESIZED_WIRE_18),
	.a4(SYNTHESIZED_WIRE_19),
	.a5(SYNTHESIZED_WIRE_20),
	.a6(SYNTHESIZED_WIRE_21),
	.a7(SYNTHESIZED_WIRE_22),
	.a8(SYNTHESIZED_WIRE_23),
	.r1(SYNTHESIZED_WIRE_24),
	.r2(SYNTHESIZED_WIRE_25),
	.r3(SYNTHESIZED_WIRE_26),
	.r4(SYNTHESIZED_WIRE_27),
	.r5(SYNTHESIZED_WIRE_28),
	.r6(SYNTHESIZED_WIRE_29),
	.r7(SYNTHESIZED_WIRE_30),
	.r8(SYNTHESIZED_WIRE_31),
	.bo_1(SYNTHESIZED_WIRE_32),
	.bo_2(SYNTHESIZED_WIRE_33),
	.bo_3(SYNTHESIZED_WIRE_34),
	.bo_4(SYNTHESIZED_WIRE_35),
	.bo_5(SYNTHESIZED_WIRE_36),
	.bo_6(SYNTHESIZED_WIRE_37),
	.bo_7(SYNTHESIZED_WIRE_38),
	.bo_8(SYNTHESIZED_WIRE_39),
	.ao_1(SYNTHESIZED_WIRE_40),
	.ao_2(SYNTHESIZED_WIRE_41),
	.ao_3(SYNTHESIZED_WIRE_42),
	.ao_4(SYNTHESIZED_WIRE_43),
	.ao_5(SYNTHESIZED_WIRE_44),
	.ao_6(SYNTHESIZED_WIRE_45),
	.ao_7(SYNTHESIZED_WIRE_46),
	.ao_8(SYNTHESIZED_WIRE_47),
	.ro_1(SYNTHESIZED_WIRE_48),
	.ro_2(SYNTHESIZED_WIRE_49),
	.ro_3(SYNTHESIZED_WIRE_50),
	.ro_4(SYNTHESIZED_WIRE_51),
	.ro_5(SYNTHESIZED_WIRE_52),
	.ro_6(SYNTHESIZED_WIRE_53),
	.ro_7(SYNTHESIZED_WIRE_54),
	.ro_8(SYNTHESIZED_WIRE_55));


multiplication_block	b2v_inst2(
	.b1(SYNTHESIZED_WIRE_32),
	.b2(SYNTHESIZED_WIRE_33),
	.b3(SYNTHESIZED_WIRE_34),
	.b4(SYNTHESIZED_WIRE_35),
	.b5(SYNTHESIZED_WIRE_36),
	.b6(SYNTHESIZED_WIRE_37),
	.b7(SYNTHESIZED_WIRE_38),
	.b8(SYNTHESIZED_WIRE_39),
	.a1(SYNTHESIZED_WIRE_40),
	.a2(SYNTHESIZED_WIRE_41),
	.a3(SYNTHESIZED_WIRE_42),
	.a4(SYNTHESIZED_WIRE_43),
	.a5(SYNTHESIZED_WIRE_44),
	.a6(SYNTHESIZED_WIRE_45),
	.a7(SYNTHESIZED_WIRE_46),
	.a8(SYNTHESIZED_WIRE_47),
	.r1(SYNTHESIZED_WIRE_48),
	.r2(SYNTHESIZED_WIRE_49),
	.r3(SYNTHESIZED_WIRE_50),
	.r4(SYNTHESIZED_WIRE_51),
	.r5(SYNTHESIZED_WIRE_52),
	.r6(SYNTHESIZED_WIRE_53),
	.r7(SYNTHESIZED_WIRE_54),
	.r8(SYNTHESIZED_WIRE_55),
	.bo_1(SYNTHESIZED_WIRE_56),
	.bo_2(SYNTHESIZED_WIRE_57),
	.bo_3(SYNTHESIZED_WIRE_58),
	.bo_4(SYNTHESIZED_WIRE_59),
	.bo_5(SYNTHESIZED_WIRE_60),
	.bo_6(SYNTHESIZED_WIRE_61),
	.bo_7(SYNTHESIZED_WIRE_62),
	.bo_8(SYNTHESIZED_WIRE_63),
	.ao_1(SYNTHESIZED_WIRE_64),
	.ao_2(SYNTHESIZED_WIRE_65),
	.ao_3(SYNTHESIZED_WIRE_66),
	.ao_4(SYNTHESIZED_WIRE_67),
	.ao_5(SYNTHESIZED_WIRE_68),
	.ao_6(SYNTHESIZED_WIRE_69),
	.ao_7(SYNTHESIZED_WIRE_70),
	.ao_8(SYNTHESIZED_WIRE_71),
	.ro_1(SYNTHESIZED_WIRE_72),
	.ro_2(SYNTHESIZED_WIRE_73),
	.ro_3(SYNTHESIZED_WIRE_74),
	.ro_4(SYNTHESIZED_WIRE_75),
	.ro_5(SYNTHESIZED_WIRE_76),
	.ro_6(SYNTHESIZED_WIRE_77),
	.ro_7(SYNTHESIZED_WIRE_78),
	.ro_8(SYNTHESIZED_WIRE_79));


multiplication_block	b2v_inst3(
	.b1(SYNTHESIZED_WIRE_56),
	.b2(SYNTHESIZED_WIRE_57),
	.b3(SYNTHESIZED_WIRE_58),
	.b4(SYNTHESIZED_WIRE_59),
	.b5(SYNTHESIZED_WIRE_60),
	.b6(SYNTHESIZED_WIRE_61),
	.b7(SYNTHESIZED_WIRE_62),
	.b8(SYNTHESIZED_WIRE_63),
	.a1(SYNTHESIZED_WIRE_64),
	.a2(SYNTHESIZED_WIRE_65),
	.a3(SYNTHESIZED_WIRE_66),
	.a4(SYNTHESIZED_WIRE_67),
	.a5(SYNTHESIZED_WIRE_68),
	.a6(SYNTHESIZED_WIRE_69),
	.a7(SYNTHESIZED_WIRE_70),
	.a8(SYNTHESIZED_WIRE_71),
	.r1(SYNTHESIZED_WIRE_72),
	.r2(SYNTHESIZED_WIRE_73),
	.r3(SYNTHESIZED_WIRE_74),
	.r4(SYNTHESIZED_WIRE_75),
	.r5(SYNTHESIZED_WIRE_76),
	.r6(SYNTHESIZED_WIRE_77),
	.r7(SYNTHESIZED_WIRE_78),
	.r8(SYNTHESIZED_WIRE_79),
	.bo_1(SYNTHESIZED_WIRE_80),
	.bo_2(SYNTHESIZED_WIRE_81),
	.bo_3(SYNTHESIZED_WIRE_82),
	.bo_4(SYNTHESIZED_WIRE_83),
	.bo_5(SYNTHESIZED_WIRE_84),
	.bo_6(SYNTHESIZED_WIRE_85),
	.bo_7(SYNTHESIZED_WIRE_86),
	.bo_8(SYNTHESIZED_WIRE_87),
	.ao_1(SYNTHESIZED_WIRE_88),
	.ao_2(SYNTHESIZED_WIRE_89),
	.ao_3(SYNTHESIZED_WIRE_90),
	.ao_4(SYNTHESIZED_WIRE_91),
	.ao_5(SYNTHESIZED_WIRE_92),
	.ao_6(SYNTHESIZED_WIRE_93),
	.ao_7(SYNTHESIZED_WIRE_94),
	.ao_8(SYNTHESIZED_WIRE_95),
	.ro_1(SYNTHESIZED_WIRE_96),
	.ro_2(SYNTHESIZED_WIRE_97),
	.ro_3(SYNTHESIZED_WIRE_98),
	.ro_4(SYNTHESIZED_WIRE_99),
	.ro_5(SYNTHESIZED_WIRE_100),
	.ro_6(SYNTHESIZED_WIRE_101),
	.ro_7(SYNTHESIZED_WIRE_102),
	.ro_8(SYNTHESIZED_WIRE_103));


multiplication_block	b2v_inst4(
	.b1(SYNTHESIZED_WIRE_80),
	.b2(SYNTHESIZED_WIRE_81),
	.b3(SYNTHESIZED_WIRE_82),
	.b4(SYNTHESIZED_WIRE_83),
	.b5(SYNTHESIZED_WIRE_84),
	.b6(SYNTHESIZED_WIRE_85),
	.b7(SYNTHESIZED_WIRE_86),
	.b8(SYNTHESIZED_WIRE_87),
	.a1(SYNTHESIZED_WIRE_88),
	.a2(SYNTHESIZED_WIRE_89),
	.a3(SYNTHESIZED_WIRE_90),
	.a4(SYNTHESIZED_WIRE_91),
	.a5(SYNTHESIZED_WIRE_92),
	.a6(SYNTHESIZED_WIRE_93),
	.a7(SYNTHESIZED_WIRE_94),
	.a8(SYNTHESIZED_WIRE_95),
	.r1(SYNTHESIZED_WIRE_96),
	.r2(SYNTHESIZED_WIRE_97),
	.r3(SYNTHESIZED_WIRE_98),
	.r4(SYNTHESIZED_WIRE_99),
	.r5(SYNTHESIZED_WIRE_100),
	.r6(SYNTHESIZED_WIRE_101),
	.r7(SYNTHESIZED_WIRE_102),
	.r8(SYNTHESIZED_WIRE_103),
	.bo_1(SYNTHESIZED_WIRE_104),
	.bo_2(SYNTHESIZED_WIRE_105),
	.bo_3(SYNTHESIZED_WIRE_106),
	.bo_4(SYNTHESIZED_WIRE_107),
	.bo_5(SYNTHESIZED_WIRE_108),
	.bo_6(SYNTHESIZED_WIRE_109),
	.bo_7(SYNTHESIZED_WIRE_110),
	.bo_8(SYNTHESIZED_WIRE_111),
	.ao_1(SYNTHESIZED_WIRE_112),
	.ao_2(SYNTHESIZED_WIRE_113),
	.ao_3(SYNTHESIZED_WIRE_114),
	.ao_4(SYNTHESIZED_WIRE_115),
	.ao_5(SYNTHESIZED_WIRE_116),
	.ao_6(SYNTHESIZED_WIRE_117),
	.ao_7(SYNTHESIZED_WIRE_118),
	.ao_8(SYNTHESIZED_WIRE_119),
	.ro_1(SYNTHESIZED_WIRE_120),
	.ro_2(SYNTHESIZED_WIRE_121),
	.ro_3(SYNTHESIZED_WIRE_122),
	.ro_4(SYNTHESIZED_WIRE_123),
	.ro_5(SYNTHESIZED_WIRE_124),
	.ro_6(SYNTHESIZED_WIRE_125),
	.ro_7(SYNTHESIZED_WIRE_126),
	.ro_8(SYNTHESIZED_WIRE_127));


multiplication_block	b2v_inst5(
	.b1(SYNTHESIZED_WIRE_104),
	.b2(SYNTHESIZED_WIRE_105),
	.b3(SYNTHESIZED_WIRE_106),
	.b4(SYNTHESIZED_WIRE_107),
	.b5(SYNTHESIZED_WIRE_108),
	.b6(SYNTHESIZED_WIRE_109),
	.b7(SYNTHESIZED_WIRE_110),
	.b8(SYNTHESIZED_WIRE_111),
	.a1(SYNTHESIZED_WIRE_112),
	.a2(SYNTHESIZED_WIRE_113),
	.a3(SYNTHESIZED_WIRE_114),
	.a4(SYNTHESIZED_WIRE_115),
	.a5(SYNTHESIZED_WIRE_116),
	.a6(SYNTHESIZED_WIRE_117),
	.a7(SYNTHESIZED_WIRE_118),
	.a8(SYNTHESIZED_WIRE_119),
	.r1(SYNTHESIZED_WIRE_120),
	.r2(SYNTHESIZED_WIRE_121),
	.r3(SYNTHESIZED_WIRE_122),
	.r4(SYNTHESIZED_WIRE_123),
	.r5(SYNTHESIZED_WIRE_124),
	.r6(SYNTHESIZED_WIRE_125),
	.r7(SYNTHESIZED_WIRE_126),
	.r8(SYNTHESIZED_WIRE_127),
	.bo_1(SYNTHESIZED_WIRE_128),
	.bo_2(SYNTHESIZED_WIRE_129),
	.bo_3(SYNTHESIZED_WIRE_130),
	.bo_4(SYNTHESIZED_WIRE_131),
	.bo_5(SYNTHESIZED_WIRE_132),
	.bo_6(SYNTHESIZED_WIRE_133),
	.bo_7(SYNTHESIZED_WIRE_134),
	.bo_8(SYNTHESIZED_WIRE_135),
	.ao_1(SYNTHESIZED_WIRE_136),
	.ao_2(SYNTHESIZED_WIRE_137),
	.ao_3(SYNTHESIZED_WIRE_138),
	.ao_4(SYNTHESIZED_WIRE_139),
	.ao_5(SYNTHESIZED_WIRE_140),
	.ao_6(SYNTHESIZED_WIRE_141),
	.ao_7(SYNTHESIZED_WIRE_142),
	.ao_8(SYNTHESIZED_WIRE_143),
	.ro_1(SYNTHESIZED_WIRE_144),
	.ro_2(SYNTHESIZED_WIRE_145),
	.ro_3(SYNTHESIZED_WIRE_146),
	.ro_4(SYNTHESIZED_WIRE_147),
	.ro_5(SYNTHESIZED_WIRE_148),
	.ro_6(SYNTHESIZED_WIRE_149),
	.ro_7(SYNTHESIZED_WIRE_150),
	.ro_8(SYNTHESIZED_WIRE_151));


multiplication_block	b2v_inst6(
	.b1(SYNTHESIZED_WIRE_128),
	.b2(SYNTHESIZED_WIRE_129),
	.b3(SYNTHESIZED_WIRE_130),
	.b4(SYNTHESIZED_WIRE_131),
	.b5(SYNTHESIZED_WIRE_132),
	.b6(SYNTHESIZED_WIRE_133),
	.b7(SYNTHESIZED_WIRE_134),
	.b8(SYNTHESIZED_WIRE_135),
	.a1(SYNTHESIZED_WIRE_136),
	.a2(SYNTHESIZED_WIRE_137),
	.a3(SYNTHESIZED_WIRE_138),
	.a4(SYNTHESIZED_WIRE_139),
	.a5(SYNTHESIZED_WIRE_140),
	.a6(SYNTHESIZED_WIRE_141),
	.a7(SYNTHESIZED_WIRE_142),
	.a8(SYNTHESIZED_WIRE_143),
	.r1(SYNTHESIZED_WIRE_144),
	.r2(SYNTHESIZED_WIRE_145),
	.r3(SYNTHESIZED_WIRE_146),
	.r4(SYNTHESIZED_WIRE_147),
	.r5(SYNTHESIZED_WIRE_148),
	.r6(SYNTHESIZED_WIRE_149),
	.r7(SYNTHESIZED_WIRE_150),
	.r8(SYNTHESIZED_WIRE_151),
	.bo_1(SYNTHESIZED_WIRE_152),
	.bo_2(SYNTHESIZED_WIRE_153),
	.bo_3(SYNTHESIZED_WIRE_154),
	.bo_4(SYNTHESIZED_WIRE_155),
	.bo_5(SYNTHESIZED_WIRE_156),
	.bo_6(SYNTHESIZED_WIRE_157),
	.bo_7(SYNTHESIZED_WIRE_158),
	.bo_8(SYNTHESIZED_WIRE_159),
	.ao_1(SYNTHESIZED_WIRE_160),
	.ao_2(SYNTHESIZED_WIRE_161),
	.ao_3(SYNTHESIZED_WIRE_162),
	.ao_4(SYNTHESIZED_WIRE_163),
	.ao_5(SYNTHESIZED_WIRE_164),
	.ao_6(SYNTHESIZED_WIRE_165),
	.ao_7(SYNTHESIZED_WIRE_166),
	.ao_8(SYNTHESIZED_WIRE_167),
	.ro_1(SYNTHESIZED_WIRE_168),
	.ro_2(SYNTHESIZED_WIRE_169),
	.ro_3(SYNTHESIZED_WIRE_170),
	.ro_4(SYNTHESIZED_WIRE_171),
	.ro_5(SYNTHESIZED_WIRE_172),
	.ro_6(SYNTHESIZED_WIRE_173),
	.ro_7(SYNTHESIZED_WIRE_174),
	.ro_8(SYNTHESIZED_WIRE_175));


multiplication_block	b2v_inst7(
	.b1(SYNTHESIZED_WIRE_152),
	.b2(SYNTHESIZED_WIRE_153),
	.b3(SYNTHESIZED_WIRE_154),
	.b4(SYNTHESIZED_WIRE_155),
	.b5(SYNTHESIZED_WIRE_156),
	.b6(SYNTHESIZED_WIRE_157),
	.b7(SYNTHESIZED_WIRE_158),
	.b8(SYNTHESIZED_WIRE_159),
	.a1(SYNTHESIZED_WIRE_160),
	.a2(SYNTHESIZED_WIRE_161),
	.a3(SYNTHESIZED_WIRE_162),
	.a4(SYNTHESIZED_WIRE_163),
	.a5(SYNTHESIZED_WIRE_164),
	.a6(SYNTHESIZED_WIRE_165),
	.a7(SYNTHESIZED_WIRE_166),
	.a8(SYNTHESIZED_WIRE_167),
	.r1(SYNTHESIZED_WIRE_168),
	.r2(SYNTHESIZED_WIRE_169),
	.r3(SYNTHESIZED_WIRE_170),
	.r4(SYNTHESIZED_WIRE_171),
	.r5(SYNTHESIZED_WIRE_172),
	.r6(SYNTHESIZED_WIRE_173),
	.r7(SYNTHESIZED_WIRE_174),
	.r8(SYNTHESIZED_WIRE_175),
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	.ro_1(r_ALTERA_SYNTHESIZED[0]),
	.ro_2(r_ALTERA_SYNTHESIZED[1]),
	.ro_3(r_ALTERA_SYNTHESIZED[2]),
	.ro_4(r_ALTERA_SYNTHESIZED[3]),
	.ro_5(r_ALTERA_SYNTHESIZED[4]),
	.ro_6(r_ALTERA_SYNTHESIZED[5]),
	.ro_7(r_ALTERA_SYNTHESIZED[6]),
	.ro_8(r_ALTERA_SYNTHESIZED[7]));


assign	r = r_ALTERA_SYNTHESIZED;

endmodule
